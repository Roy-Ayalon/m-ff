//-----------------------------------------------------------------------------
// Project       : Register Test Bench
//-----------------------------------------------------------------------------
// File          : register_test_bench.v
// Author        : Roy Ayalon 
// Created       : 23 March 2023
//-----------------------------------------------------------------------------

module tb;  

// -----------------------------------------------------------------------------
// Parameter / Define
// -----------------------------------------------------------------------------

parameter       WIDTH = 12;         //Width of data path
parameter       RESET_VAL = 0;      //Reset value for data path

// -----------------------------------------------------------------------------
// Register/Wires Declarations
// -----------------------------------------------------------------------------

reg                             clk;
reg                             rst_n;
reg                             enable;
reg  [WIDTH-1:0]                data_in;

wire [WIDTH-1:0]                data_out;

// -----------------------------------------------------------------------------
// clock / reset generator
// -----------------------------------------------------------------------------

always #5 clk = ~clk;

// -----------------------------------------------------------------------------
//  DUT
// -----------------------------------------------------------------------------

m_ff #(.WIDTH(WIDTH), .RESET_VAL(RESET_VAL)) m_ff (
.clk(clk),
.rst_n(rst_n),
.enable(enable),
.data_in(data_in),
.data_out(data_out));

// -----------------------------------------------------------------------------
//  Sim Base Run
// -----------------------------------------------------------------------------

initial begin
$display("TEST STARTED");
clk = 0;
rst_n = 0;
enable = 0;
data_in = 0;


repeat (5) @(posedge clk);
#1;
rst_n = 1;

repeat (5) @(posedge clk);
data_in =#1 750;
repeat (7) @(posedge clk);
data_in =#1 302;
enable = 1;

repeat (7) @(posedge clk);
$display("TEST FINISHED");
$finish;
end

// -----------------------------------------------------------------------------
//  Waves
// -----------------------------------------------------------------------------
initial begin
$dumpfile("tb.vcd");
$dumpvars(1,tb);
end 


// -----------------------------------------------------------------------------
//  Checkers
// -----------------------------------------------------------------------------

// -----------------------------------------------------------------------------
//  TASKS & Functions
// -----------------------------------------------------------------------------



endmodule

